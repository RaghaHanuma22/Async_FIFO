#module for synchronizer
