#Module for write pointerr
