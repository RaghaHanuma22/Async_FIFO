#module for read pointer
