#Module for fifo memory
#Author: Raghav
