#Testbench - Conventional for sanity check
