`include "uvm_macros.svh"
import uvm_pkg::*;

package rd_pkg;
    `include "rd_seq_item.sv"
    `include "rd_sequence.sv"
    `include "rd_monitor.sv"
    `include "rd_driver.sv"
    `include "rd_agent.sv"
endpackage

