#Top module
